// Ps2.v

// Generated using ACDS version 23.1 993

`timescale 1 ps / 1 ps
module Ps2 (
		input  wire [7:0] command,       // avalon_ps2_command_sink.data
		input  wire       command_valid, //                        .valid
		output wire       command_ready, //                        .ready
		input  wire       data_ready,    //  avalon_ps2_data_source.ready
		output wire [7:0] data,          //                        .data
		output wire       data_valid,    //                        .valid
		input  wire       clk,           //                     clk.clk
		inout  wire       PS2_CLK,       //      external_interface.CLK
		inout  wire       PS2_DAT,       //                        .DAT
		input  wire       reset          //                   reset.reset
	);

	Ps2_ps2_0 ps2_0 (
		.clk           (clk),           //                     clk.clk
		.reset         (reset),         //                   reset.reset
		.command       (command),       // avalon_ps2_command_sink.data
		.command_valid (command_valid), //                        .valid
		.command_ready (command_ready), //                        .ready
		.data_ready    (data_ready),    //  avalon_ps2_data_source.ready
		.data          (data),          //                        .data
		.data_valid    (data_valid),    //                        .valid
		.PS2_CLK       (PS2_CLK),       //      external_interface.export
		.PS2_DAT       (PS2_DAT)        //                        .export
	);

endmodule
